module iic_tx (

);

endmodule : iic_tx
