`timescale 1ns / 1ps

module AimBot (
);

endmodule : AimBot
