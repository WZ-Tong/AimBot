module GTP_IOCLKBUF #(parameter GATE_EN = "FALSE") (
    output CLKOUT,
    input  CLKIN ,
    input  DI
);

endmodule : GTP_IOCLKBUF
