module GTP_OUTBUFT (
    output O,
    input I,
    input T
);
    parameter IOSTANDARD = "DEFAULT";
    parameter SLEW_RATE = "SLOW";
    parameter DRIVE_STRENGTH = "8";
endmodule
