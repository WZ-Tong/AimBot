module pll (
    input  clkin1  ,
    input  pll_rst ,

    output pll_lock,
    output clkout0 ,
    output clkout1
);

endmodule : pll
