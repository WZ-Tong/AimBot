module GTP_INBUF (
    output O,
    input I
);
    parameter IOSTANDARD = "DEFAULT";
    parameter TERM_DDR = "ON";
endmodule
