module GTP_IOCLKDIV #(
    parameter GRS_EN     = "TRUE",
    parameter DIV_FACTOR = "2"
) (
    output CLKDIVOUT,
    input  CLKIN    ,
    input  RST_N
);

endmodule : GTP_IOCLKDIV
