module GTP_INBUFG (
    output O,
    input I
);
    parameter IOSTANDARD = "DEFAULT";
    parameter TERM_DDR = "ON";
endmodule
