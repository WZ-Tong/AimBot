module GTP_CLKBUFG (
    output CLKOUT,
    input CLKIN
);
endmodule
