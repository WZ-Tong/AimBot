module ddr3 #(
    parameter  DATA_WIDTH = 16                                               ,
    localparam DM_WIDTH   = DATA_WIDTH==16 ? 2 : (DATA_WIDTH==32 ? 4 : 0)    ,
    localparam DQ_WIDTH   = DATA_WIDTH==16 ? 2 : (DATA_WIDTH==32 ? 4 : 0)    ,
    localparam DATA_LEN   = DATA_WIDTH==16 ? 128 : (DATA_WIDTH==32 ? 256 : 0)
) (
    input                   clk            ,
    output                  inited         ,
    output                  phy_clk        ,
    output                  phy_clkl       ,

    input  [          27:0] axi_awaddr     ,
    input  [           3:0] axi_awlen      ,
    output                  axi_awready    ,
    input                   axi_awvalid    ,

    input  [  DATA_LEN-1:0] axi_wdata      ,
    input  [DATA_WIDTH-1:0] axi_wstrb      ,
    output                  axi_wready     ,
    output                  axi_wusero_last,

    input  [          27:0] axi_araddr     ,
    input  [           3:0] axi_arlen      ,
    output                  axi_arready    ,
    input                   axi_arvalid    ,

    output [  DATA_LEN-1:0] axi_rdata      ,
    output [           3:0] axi_rid        ,
    output                  axi_rlast      ,
    output                  axi_rvalid     ,

    output                  mem_rst_n      ,
    output                  mem_ck         ,
    output                  mem_ck_n       ,
    output                  mem_cke        ,
    output                  mem_cs_n       ,
    output                  mem_ras_n      ,
    output                  mem_cas_n      ,
    output                  mem_we_n       ,
    output                  mem_odt        ,

    output [          14:0] mem_a          ,
    output [           2:0] mem_ba         ,
    inout  [  DQ_WIDTH-1:0] mem_dqs        ,
    inout  [  DQ_WIDTH-1:0] mem_dqs_n      ,
    inout  [DATA_WIDTH-1:0] mem_dq         ,
    output [  DM_WIDTH-1:0] mem_dm
);

    if (DATA_WIDTH==16) begin : gen_ddr3_16
        ddr3_16 u_ddr3_16 (
            .clk            (clk            ),
            .inited         (inited         ),
            .phy_clk        (phy_clk        ),
            .phy_clkl       (phy_clkl       ),
            .axi_awaddr     (axi_awaddr     ),
            .axi_awlen      (axi_awlen      ),
            .axi_awready    (axi_awready    ),
            .axi_awvalid    (axi_awvalid    ),
            .axi_wdata      (axi_wdata      ),
            .axi_wstrb      (axi_wstrb      ),
            .axi_wready     (axi_wready     ),
            .axi_wusero_last(axi_wusero_last),
            .axi_araddr     (axi_araddr     ),
            .axi_arlen      (axi_arlen      ),
            .axi_arready    (axi_arready    ),
            .axi_arvalid    (axi_arvalid    ),
            .axi_rdata      (axi_rdata      ),
            .axi_rid        (axi_rid        ),
            .axi_rlast      (axi_rlast      ),
            .axi_rvalid     (axi_rvalid     ),
            .mem_rst_n      (mem_rst_n      ),
            .mem_ck         (mem_ck         ),
            .mem_ck_n       (mem_ck_n       ),
            .mem_cke        (mem_cke        ),
            .mem_cs_n       (mem_cs_n       ),
            .mem_ras_n      (mem_ras_n      ),
            .mem_cas_n      (mem_cas_n      ),
            .mem_we_n       (mem_we_n       ),
            .mem_odt        (mem_odt        ),
            .mem_a          (mem_a          ),
            .mem_ba         (mem_ba         ),
            .mem_dqs        (mem_dqs        ),
            .mem_dqs_n      (mem_dqs_n      ),
            .mem_dq         (mem_dq         ),
            .mem_dm         (mem_dm         )
        );
    end else if (DATA_WIDTH==32) begin : gen_ddr3_32
        ddr3_32 u_ddr3_32 (
            .clk            (clk            ),
            .inited         (inited         ),
            .phy_clk        (phy_clk        ),
            .phy_clkl       (phy_clkl       ),
            .axi_awaddr     (axi_awaddr     ),
            .axi_awlen      (axi_awlen      ),
            .axi_awready    (axi_awready    ),
            .axi_awvalid    (axi_awvalid    ),
            .axi_wdata      (axi_wdata      ),
            .axi_wstrb      (axi_wstrb      ),
            .axi_wready     (axi_wready     ),
            .axi_wusero_last(axi_wusero_last),
            .axi_araddr     (axi_araddr     ),
            .axi_arlen      (axi_arlen      ),
            .axi_arready    (axi_arready    ),
            .axi_arvalid    (axi_arvalid    ),
            .axi_rdata      (axi_rdata      ),
            .axi_rid        (axi_rid        ),
            .axi_rlast      (axi_rlast      ),
            .axi_rvalid     (axi_rvalid     ),
            .mem_rst_n      (mem_rst_n      ),
            .mem_ck         (mem_ck         ),
            .mem_ck_n       (mem_ck_n       ),
            .mem_cke        (mem_cke        ),
            .mem_cs_n       (mem_cs_n       ),
            .mem_ras_n      (mem_ras_n      ),
            .mem_cas_n      (mem_cas_n      ),
            .mem_we_n       (mem_we_n       ),
            .mem_odt        (mem_odt        ),
            .mem_a          (mem_a          ),
            .mem_ba         (mem_ba         ),
            .mem_dqs        (mem_dqs        ),
            .mem_dqs_n      (mem_dqs_n      ),
            .mem_dq         (mem_dq         ),
            .mem_dm         (mem_dm         )
        );
    end

endmodule : ddr3
