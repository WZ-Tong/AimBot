module AimBot (
);

endmodule : AimBot
