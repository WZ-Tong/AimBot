module pll (
    input  clkin1  ,
    input  pll_rst ,

    output pll_lock,
    output clkout0 ,
    output clkout1 ,
    output clkout2
);

endmodule : pll
