module rgmii_stat (
    input  clk   ,
    input  inited,
    input  error ,
    input  tx    ,
    input  rx    ,

    output stat
);

endmodule : rgmii_stat
